module cam_decorder#()();



endmodule // cam_decorder
