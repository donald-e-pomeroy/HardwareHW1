module flipflop(data_i, data_o);
   


  
  endmodule; // flipflop




