module cam(read_i, 
	   read_index_i, 
	   write_i, 
	   write_index_i, 
	   write_data_i, 
	   search_i, 
	   search_data_i, 
	   read_valid_o,
	   read_value_o,
	   search_valid_o
	   search_index_o);

   

  endmodule