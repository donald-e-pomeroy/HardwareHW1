module cam()

  endmodule