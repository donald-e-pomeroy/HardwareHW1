module flipflop()

  endmodule; // flipflop




