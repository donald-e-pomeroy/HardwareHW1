module flipflop()

  endmodule; // flipflop


